module and1(dataIn1, dataIn2, dataOut);
input dataIn1, dataIn2;
output dataOut;
assign dataOut = dataIn1 & dataIn2;
endmodule
